module and1(i1,i2,saida);
input i1, i2;
output saida;
assign saida=(i1&i2)?1:0;




endmodule // and
